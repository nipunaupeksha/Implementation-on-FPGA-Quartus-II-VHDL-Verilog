library ieee;
use ieee.std_logic_1164.all;
entity prio_encoder42 is
    port(r:in std_logic_vector(3 downto 0);
    code: out std_logic_vector(1 downto 0);
    active: out std_logic);
    end prio_encoder42;

    architecture cond_arch of prio_encoder42 is
        begin
            code<="11" when (r(3)='1') else
                "10" when (r(2)='1') else
                "00" when (r(1)='1') else
                "00";
            active<=r(3) or r(2) or r(1) or r(0);
            end cond_arch;
